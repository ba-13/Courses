// Hello world to verilog

module hello ();

  initial
    $display("Hello Verilog!");

endmodule

