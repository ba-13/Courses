module feed_forward (A, B);
    input A;
    output B;
    assign B = A;
endmodule